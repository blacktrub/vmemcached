module vmemcached

import net

pub struct Connection {
	host string = '127.0.0.1'
	port int = 11211
}

pub struct Memcached {
	socket net.Socket
}

pub struct Value {
pub:
	content string
}

fn clean_response(response string) string {
	return response.replace('\r\n', '')
}

pub fn connect(opt Connection) ?Memcached {
	socket := net.dial(opt.host, opt.port) or {
		return error(err)
	}
	return Memcached{
		socket: socket
	}
}

pub fn (m Memcached) disconnect() {
	m.socket.close() or { }
}

pub fn (m Memcached) flushall() bool {
	message := 'flush_all\r\n'
	m.socket.write(message) or {
		return false
	}
	response := m.socket.read_line()[0..2]
	return match response {
		'OK' { true }
		else { false }
	}
}

pub fn (m Memcached) get(key string) Value {
	msg := 'get $key\r\n'
	m.socket.write(msg) or {
		return Value{}
	}
	response := m.socket.read_line()
	if response == 'END\r\n' {
		return Value{}
	}
	// TODO: why?
	m.socket.read_line()
	value := m.socket.read_line()
	return Value{clean_response(value)}
}

pub fn (m Memcached) set(key, val string) bool {
	msg := 'set $key 0 0 $val.len\r\n$val\r\n'
	m.socket.write(msg) or {
		return false
	}
	response := m.socket.read_line()[0..6]
	return match response {
		'STORED' { true }
		else { false }
	}
}

pub fn (m Memcached) replace(key, val string) bool {
	msg := 'replace $key 0 0 $val.len\r\n$val\r\n'
	m.socket.write(msg) or {
		return false
	}
	// TODO: why?
	// see https://github.com/vlang/v/blob/master/vlib/net/socket.v#L310
	m.socket.read_line()
	response := clean_response(m.socket.read_line())
	return match response {
		'STORED' { true }
		else { false }
	}
}

pub fn (m Memcached) delete(key string) bool {
	msg := 'delete $key\r\n'
	m.socket.write(msg) or {
		return false
	}
	m.socket.read_line()
	response := clean_response(m.socket.read_line())
	return match response {
		'DELETED' { true }
		else { false }
	}
}

pub fn (m Memcached) add(key, val string) bool {
	msg := 'add $key 0 0 $val.len\r\n$val'
	m.socket.write(msg) or {
		return false
	}
	response := clean_response(m.socket.read_line())
	return match response {
		'STORED' { true }
		else { false }
	}
}

pub fn (m Memcached) incr(key, val string) bool {
	msg := 'incr $key $val'
	m.socket.write(msg) or {
		return false
	}
	response := clean_response(m.socket.read_line())
	return match response {
		'NOT_FOUND' { false }
		else { true }
	}
}

pub fn (m Memcached) decr(key, val string) bool {
	msg := 'decr $key $val'
	m.socket.write(msg) or {
		return false
	}
	response := clean_response(m.socket.read_line())
	return match response {
		'NOT_FOUND' { false }
		else { true }
	}
}
